-- r-VEX processor MMU
-- Copyright (C) 2008-2016 by TU Delft.
-- All Rights Reserved.

-- THIS IS A LEGAL DOCUMENT, BY USING r-VEX,
-- YOU ARE AGREEING TO THESE TERMS AND CONDITIONS.

-- No portion of this work may be used by any commercial entity, or for any
-- commercial purpose, without the prior, written permission of TU Delft.
-- Nonprofit and noncommercial use is permitted as described below.

-- 1. r-VEX is provided AS IS, with no warranty of any kind, express
-- or implied. The user of the code accepts full responsibility for the
-- application of the code and the use of any results.

-- 2. Nonprofit and noncommercial use is encouraged. r-VEX may be
-- downloaded, compiled, synthesized, copied, and modified solely for nonprofit,
-- educational, noncommercial research, and noncommercial scholarship
-- purposes provided that this notice in its entirety accompanies all copies.
-- Copies of the modified software can be delivered to persons who use it
-- solely for nonprofit, educational, noncommercial research, and
-- noncommercial scholarship purposes provided that this notice in its
-- entirety accompanies all copies.

-- 3. ALL COMMERCIAL USE, AND ALL USE BY FOR PROFIT ENTITIES, IS EXPRESSLY
-- PROHIBITED WITHOUT A LICENSE FROM TU Delft (J.S.S.M.Wong@tudelft.nl).

-- 4. No nonprofit user may place any restrictions on the use of this software,
-- including as modified by the user, by any other authorized user.

-- 5. Noncommercial and nonprofit users may distribute copies of r-VEX
-- in compiled or binary form as set forth in Section 2, provided that
-- either: (A) it is accompanied by the corresponding machine-readable source
-- code, or (B) it is accompanied by a written offer, with no time limit, to
-- give anyone a machine-readable copy of the corresponding source code in
-- return for reimbursement of the cost of distribution. This written offer
-- must permit verbatim duplication by anyone, or (C) it is distributed by
-- someone who received only the executable form, and is accompanied by a
-- copy of the written offer of source code.

-- 6. r-VEX was developed by Stephan Wong, Thijs van As, Fakhar Anjam,
-- Roel Seedorf, Anthony Brandon, Jeroen van Straten. r-VEX is currently
-- maintained by TU Delft (J.S.S.M.Wong@tudelft.nl).

-- 7. The MMU was created by Jens Johansen.

-- Copyright (C) 2008-2016 by TU Delft.

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library rvex;
use rvex.cache_pkg.all;

--=============================================================================
-- This entity represents a content-addressable memory, used by the CAM. It is
-- implemented using block RAMs. A 10-bit input (data) and a 5-bit output
-- (address) results in one block RAM. Essentially, the data is used as the
-- address of the block RAM, and the associated address is one-hot encoded in
-- the block RAM data. When the data needs to be larger than 10 bits, the
-- data is split into multiple parts, each fed to a different block RAM.
-- Because the indices are one-hot encoded, the block RAM outputs can just be
-- ANDed together. This results in linear resource utilization versus data
-- width instead of exponential. The address is returned still in one-hot
-- format, to allow multiple CAMs to work together. This allows some of those
-- individual CAMs to be conditionally ignored.
-------------------------------------------------------------------------------
entity cache_tlb_cam is
--=============================================================================
  generic (
    
    -- Width of the data that is to be looked up.
    DATA_WIDTH                  : natural := 10;
    
    -- Width of the address in bits = the log2 of the number of entries.
    ADDRESS_WIDTH               : natural := 5
    
  );
  port (
    
    ---------------------------------------------------------------------------
    -- System control
    ---------------------------------------------------------------------------
    -- Active high synchronous reset input.
    reset                       : in  std_logic;
    
    -- Clock input, registers are rising edge triggered.
    clk                         : in  std_logic;
    
    -- Active high global clock enable input.
    clkEn                       : in  std_logic;
    
    ---------------------------------------------------------------------------
    -- CAM ports
    ---------------------------------------------------------------------------
    -- Data input for lookup and modification.
    data                        : in  std_logic_vector(DATA_WIDTH-1 downto 0);
    
    -- One-hot encoded address output, valid one clkEn'd cycle after data.
    addr                        : out std_logic_vector(2**ADDRESS_WIDTH-1 downto 0)
    
    -- TODO

  );
end cache_tlb_cam;

--=============================================================================
architecture arch of cache_tlb_cam is
--=============================================================================


--=============================================================================
begin -- architecture
--=============================================================================
  

end architecture;
