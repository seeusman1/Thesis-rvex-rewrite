library IEEE;
use IEEE.std_logic_1164.all;

package tta0_gcu_opcodes is
  constant IFE_CALL : integer := 0;
  constant IFE_JUMP : integer := 1;
end tta0_gcu_opcodes;
