../../lib/rvex/core/core_pipeline_pkg.template.vhd