../../lib/rvex/core/core_ctrlRegs_pkg.template.vhd