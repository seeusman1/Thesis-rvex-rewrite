-- r-VEX processor
-- Copyright (C) 2008-2014 by TU Delft.
-- All Rights Reserved.

-- THIS IS A LEGAL DOCUMENT, BY USING r-VEX,
-- YOU ARE AGREEING TO THESE TERMS AND CONDITIONS.

-- No portion of this work may be used by any commercial entity, or for any
-- commercial purpose, without the prior, written permission of TU Delft.
-- Nonprofit and noncommercial use is permitted as described below.

-- 1. r-VEX is provided AS IS, with no warranty of any kind, express
-- or implied. The user of the code accepts full responsibility for the
-- application of the code and the use of any results.

-- 2. Nonprofit and noncommercial use is encouraged. r-VEX may be
-- downloaded, compiled, synthesized, copied, and modified solely for nonprofit,
-- educational, noncommercial research, and noncommercial scholarship
-- purposes provided that this notice in its entirety accompanies all copies.
-- Copies of the modified software can be delivered to persons who use it
-- solely for nonprofit, educational, noncommercial research, and
-- noncommercial scholarship purposes provided that this notice in its
-- entirety accompanies all copies.

-- 3. ALL COMMERCIAL USE, AND ALL USE BY FOR PROFIT ENTITIES, IS EXPRESSLY
-- PROHIBITED WITHOUT A LICENSE FROM TU Delft (J.S.S.M.Wong@tudelft.nl).

-- 4. No nonprofit user may place any restrictions on the use of this software,
-- including as modified by the user, by any other authorized user.

-- 5. Noncommercial and nonprofit users may distribute copies of r-VEX
-- in compiled or binary form as set forth in Section 2, provided that
-- either: (A) it is accompanied by the corresponding machine-readable source
-- code, or (B) it is accompanied by a written offer, with no time limit, to
-- give anyone a machine-readable copy of the corresponding source code in
-- return for reimbursement of the cost of distribution. This written offer
-- must permit verbatim duplication by anyone, or (C) it is distributed by
-- someone who received only the executable form, and is accompanied by a
-- copy of the written offer of source code.

-- 6. r-VEX was developed by Stephan Wong, Thijs van As, Fakhar Anjam,
-- Roel Seedorf, Anthony Brandon, Jeroen van Straten. r-VEX is currently
-- maintained by TU Delft (J.S.S.M.Wong@tudelft.nl).

-- Copyright (C) 2008-2014 by TU Delft.

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;

library rvex;
use rvex.bus_pkg.all;

--=============================================================================
-- This peripheral provides a debugging interface between one or more rvex
-- processors and a computer, utilizing a (by default) 115200 baud UART. The
-- application(s) running on the processor can send and receive bytes to and
-- from this unit as if it were a normal UART with FIFO and interrupts, but the
-- computer can also send debugging requests and receive replies over the same
-- link. These requests and replies are handled and generated by hardware - the
-- application does not need to be aware of the existence of these packets. The
-- packets are marked in the bytestream using unique control characters; when
-- the application desires to send one of these characters, they are
-- appropriately escaped in hardware.
-------------------------------------------------------------------------------
entity periph_uart is
--=============================================================================
  generic (
    
    -- Input clock frequency.
    F_CLK                       : real := 75000000.0;
    
    -- Desired baud rate. The input clock frequency must be at least 8 times as
    -- high.
    F_BAUD                      : real := 115200.0
    
  );
  port (
    
    ---------------------------------------------------------------------------
    -- System control
    ---------------------------------------------------------------------------
    -- Active high synchronous reset input.
    reset                       : in  std_logic;
    
    -- Clock input, registers are rising edge triggered.
    clk                         : in  std_logic;
    
    -- Active high global clock enable input.
    clkEn                       : in  std_logic;
    
    ---------------------------------------------------------------------------
    -- UART pins
    ---------------------------------------------------------------------------
    -- Receive data.
    rx                          : in  std_logic;
    
    -- Transmit data.
    tx                          : out std_logic;
    
    ---------------------------------------------------------------------------
    -- Slave bus
    ---------------------------------------------------------------------------
    -- The UART can be accessed from this bus for transmitting user data over
    -- the same physical line as the debug data. Refer to the entity
    -- description in periph_uart_busIface.vhd for more information.
    -- Slave bus port.
    bus2uart                    : in  bus_mst2slv_type;
    uart2bus                    : out bus_slv2mst_type;
    
    -- Active high interrupt request output.
    irq                         : out std_logic;
    
    ---------------------------------------------------------------------------
    -- Debug interface
    ---------------------------------------------------------------------------
    -- This bus master is controlled by the debug packets, to allow the
    -- debugging software running on the computer to access mapped memory
    -- regions.
    uart2dbg_bus                : out bus_mst2slv_type;
    dbg2uart_bus                : in  bus_slv2mst_type
    
  );
end periph_uart;

--=============================================================================
architecture Behavioral of periph_uart is
--=============================================================================
  
  -- UART <-> switch signals.
  signal uart2sw_rxData         : std_logic_vector(7 downto 0);
  signal uart2sw_rxFrameError   : std_logic;
  signal uart2sw_rxStrobe       : std_logic;
  signal sw2uart_txData         : std_logic_vector(7 downto 0);
  signal sw2uart_txStrobe       : std_logic;
  signal uart2sw_txBusy         : std_logic;
  
  -- Switch/UART <-> bus interface signals.
  signal sw2user_rxData         : std_logic_vector(7 downto 0);
  signal sw2user_rxStrobe       : std_logic;
  signal user2sw_txData         : std_logic_vector(7 downto 0);
  signal user2sw_txStrobe       : std_logic;
  signal sw2user_txBusy         : std_logic;
  signal uart2user_rxCharTimeout: std_logic;
  
  -- Switch <-> debug packet controller signals.
  signal sw2pkctrl_rxData       : std_logic_vector(7 downto 0);
  signal sw2pkctrl_rxEndPacket  : std_logic;
  signal sw2pkctrl_rxStrobe     : std_logic;
  signal pkctrl2sw_txData       : std_logic_vector(7 downto 0);
  signal pkctrl2sw_txStartPacket: std_logic;
  signal pkctrl2sw_txRequest    : std_logic;
  signal sw2pkctrl_txAck        : std_logic;
  
  -- Debug packet controller <-> debug packet handler signals.
  signal pkctrl2pkhan_rxData    : std_logic_vector(7 downto 0);
  signal pkhan2pkctrl_rxPop     : std_logic;
  signal pkctrl2pkhan_rxEmpty   : std_logic;
  signal pkctrl2pkhan_rxSwap    : std_logic;
  signal pkhan2pkctrl_rxReady   : std_logic;
  signal pkhan2pkctrl_txData    : std_logic_vector(7 downto 0);
  signal pkhan2pkctrl_txPush    : std_logic;
  signal pkctrl2pkhan_txFull    : std_logic;
  signal pkctrl2pkhan_txReset   : std_logic;
  signal pkctrl2pkhan_txSwap    : std_logic;
  signal pkhan2pkctrl_txReady   : std_logic;
  
--=============================================================================
begin -- architecture
--=============================================================================
  
  -----------------------------------------------------------------------------
  -- Instantiate the UART
  -----------------------------------------------------------------------------
  uart_inst: entity rvex.utils_uart
    generic map (
      F_CLK                     => F_CLK,
      F_BAUD                    => F_BAUD,
      ENABLE_TX                 => true,
      ENABLE_RX                 => true
    )
    port map (
      
      -- System control.
      reset                     => reset,
      clk                       => clk,
      clkEn                     => clkEn,
      
      -- External interface.
      rx                        => rx,
      tx                        => tx,
      
      -- RX logic internal interface.
      rx_data                   => uart2sw_rxData,
      rx_frameError             => uart2sw_rxFrameError,
      rx_strobe                 => uart2sw_rxStrobe,
      rx_charTimeout            => uart2user_rxCharTimeout,
      
      -- TX logic internal interface.
      tx_data                   => sw2uart_txData,
      tx_strobe                 => sw2uart_txStrobe,
      tx_busy                   => uart2sw_txBusy
      
    );
  
  -----------------------------------------------------------------------------
  -- Instantiate the bytestream switch
  -----------------------------------------------------------------------------
  -- This inserts and handles special control characters and escape sequences
  -- for them to switch between transmitting/receicing application data and
  -- debug packets.
  uart_switch_inst: entity rvex.periph_uart_switch
    port map (
      
      -- System control.
      reset                     => reset,
      clk                       => clk,
      clkEn                     => clkEn,
      
      -- RX interface.
      uart2sw_rxData            => uart2sw_rxData,
      uart2sw_rxFrameError      => uart2sw_rxFrameError,
      uart2sw_rxStrobe          => uart2sw_rxStrobe,
      
      sw2user_rxData            => sw2user_rxData,
      sw2user_rxStrobe          => sw2user_rxStrobe,
      
      sw2dbg_rxData             => sw2pkctrl_rxData,
      sw2dbg_rxEndPacket        => sw2pkctrl_rxEndPacket,
      sw2dbg_rxStrobe           => sw2pkctrl_rxStrobe,
      
      -- TX interface.
      sw2uart_txData            => sw2uart_txData,
      sw2uart_txStrobe          => sw2uart_txStrobe,
      uart2sw_txBusy            => uart2sw_txBusy,
      
      user2sw_txData            => user2sw_txData,
      user2sw_txStrobe          => user2sw_txStrobe,
      sw2user_txBusy            => sw2user_txBusy,
      
      dbg2sw_txData             => pkctrl2sw_txData,
      dbg2sw_txStartPacket      => pkctrl2sw_txStartPacket,
      dbg2sw_txRequest          => pkctrl2sw_txRequest,
      sw2dbg_txAck              => sw2pkctrl_txAck
      
    );
  
  -----------------------------------------------------------------------------
  -- Instantiate the debug packet controller
  -----------------------------------------------------------------------------
  -- This handles CRC generation/verification and buffering of debug packets.
  debug_packet_control_inst: entity rvex.periph_uart_packetControl
    port map (
      
      -- System control.
      reset                     => reset,
      clk                       => clk,
      clkEn                     => clkEn,
      
      -- Interface with the packet handler.
      pkctrl2pkhan_rxData       => pkctrl2pkhan_rxData,
      pkhan2pkctrl_rxPop        => pkhan2pkctrl_rxPop,
      pkctrl2pkhan_rxEmpty      => pkctrl2pkhan_rxEmpty,
      pkctrl2pkhan_rxSwap       => pkctrl2pkhan_rxSwap,
      pkhan2pkctrl_rxReady      => pkhan2pkctrl_rxReady,
      pkhan2pkctrl_txData       => pkhan2pkctrl_txData,
      pkhan2pkctrl_txPush       => pkhan2pkctrl_txPush,
      pkctrl2pkhan_txFull       => pkctrl2pkhan_txFull,
      pkctrl2pkhan_txReset      => pkctrl2pkhan_txReset,
      pkctrl2pkhan_txSwap       => pkctrl2pkhan_txSwap,
      pkhan2pkctrl_txReady      => pkhan2pkctrl_txReady,
      
      -- Interface with UART stream switch.
      sw2pkctrl_rxData          => sw2pkctrl_rxData,
      sw2pkctrl_rxEndPacket     => sw2pkctrl_rxEndPacket,
      sw2pkctrl_rxStrobe        => sw2pkctrl_rxStrobe,
      pkctrl2sw_txData          => pkctrl2sw_txData,
      pkctrl2sw_txStartPacket   => pkctrl2sw_txStartPacket,
      pkctrl2sw_txRequest       => pkctrl2sw_txRequest,
      sw2pkctrl_txAck           => sw2pkctrl_txAck
      
    );
  
  -----------------------------------------------------------------------------
  -- Instantiate the debug packet handler
  -----------------------------------------------------------------------------
  -- This converts the incoming debug packets into bus accesses.
  debug_packet_handler: entity rvex.periph_uart_packetHandler
    port map (
      
      -- System control.
      reset                     => reset,
      clk                       => clk,
      clkEn                     => clkEn,
      
      -- Interface with packet control.
      pkctrl2pkhan_rxData       => pkctrl2pkhan_rxData,
      pkhan2pkctrl_rxPop        => pkhan2pkctrl_rxPop,
      pkctrl2pkhan_rxEmpty      => pkctrl2pkhan_rxEmpty,
      pkctrl2pkhan_rxSwap       => pkctrl2pkhan_rxSwap,
      pkhan2pkctrl_rxReady      => pkhan2pkctrl_rxReady,
      pkhan2pkctrl_txData       => pkhan2pkctrl_txData,
      pkhan2pkctrl_txPush       => pkhan2pkctrl_txPush,
      pkctrl2pkhan_txFull       => pkctrl2pkhan_txFull,
      pkctrl2pkhan_txReset      => pkctrl2pkhan_txReset,
      pkctrl2pkhan_txSwap       => pkctrl2pkhan_txSwap,
      pkhan2pkctrl_txReady      => pkhan2pkctrl_txReady,
      
      -- Bus interface.
      pkhan2dbg_bus             => uart2dbg_bus,
      dbg2pkhan_bus             => dbg2uart_bus
      
    );
  
  -----------------------------------------------------------------------------
  -- Instantiate the bus interface
  -----------------------------------------------------------------------------
  -- This will interface between the slave bus interface which the application
  -- can access to transmit and receive bytes, and the UART stream switch.
  bus_interface: entity rvex.periph_uart_busIface
    port map (
      
      -- System control.
      reset                     => reset,
      clk                       => clk,
      clkEn                     => clkEn,
      
      -- Slave bus.
      bus2uart                  => bus2uart,
      uart2bus                  => uart2bus,
      irq                       => irq,
      
      -- UART data inferface.
      rxData                    => sw2user_rxData,
      rxStrobe                  => sw2user_rxStrobe,
      rxTimeout                 => uart2user_rxCharTimeout,
      txData                    => user2sw_txData,
      txStrobe                  => user2sw_txStrobe,
      txBusy                    => sw2user_txBusy
      
    );
  
end Behavioral;
