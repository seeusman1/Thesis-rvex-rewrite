../../lib/rvex/core/core_globalRegLogic.template.vhd