package tta0_params is
  constant fu_LSU_dataw : integer := 32;
  constant fu_LSU_addrw : integer := 15;
  constant fu_stdout_dataw : integer := 8;
  constant fu_stdout_addrw : integer := 10;
  constant fu_LSU_PARAM_dataw : integer := 32;
  constant fu_LSU_PARAM_addrw : integer := 11;
end tta0_params;
