../../lib/rvex/core/core_trap_pkg.template.vhd