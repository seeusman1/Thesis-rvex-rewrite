-- r-VEX processor MMU
-- Copyright (C) 2008-2016 by TU Delft.
-- All Rights Reserved.

-- THIS IS A LEGAL DOCUMENT, BY USING r-VEX,
-- YOU ARE AGREEING TO THESE TERMS AND CONDITIONS.

-- No portion of this work may be used by any commercial entity, or for any
-- commercial purpose, without the prior, written permission of TU Delft.
-- Nonprofit and noncommercial use is permitted as described below.

-- 1. r-VEX is provided AS IS, with no warranty of any kind, express
-- or implied. The user of the code accepts full responsibility for the
-- application of the code and the use of any results.

-- 2. Nonprofit and noncommercial use is encouraged. r-VEX may be
-- downloaded, compiled, synthesized, copied, and modified solely for nonprofit,
-- educational, noncommercial research, and noncommercial scholarship
-- purposes provided that this notice in its entirety accompanies all copies.
-- Copies of the modified software can be delivered to persons who use it
-- solely for nonprofit, educational, noncommercial research, and
-- noncommercial scholarship purposes provided that this notice in its
-- entirety accompanies all copies.

-- 3. ALL COMMERCIAL USE, AND ALL USE BY FOR PROFIT ENTITIES, IS EXPRESSLY
-- PROHIBITED WITHOUT A LICENSE FROM TU Delft (J.S.S.M.Wong@tudelft.nl).

-- 4. No nonprofit user may place any restrictions on the use of this software,
-- including as modified by the user, by any other authorized user.

-- 5. Noncommercial and nonprofit users may distribute copies of r-VEX
-- in compiled or binary form as set forth in Section 2, provided that
-- either: (A) it is accompanied by the corresponding machine-readable source
-- code, or (B) it is accompanied by a written offer, with no time limit, to
-- give anyone a machine-readable copy of the corresponding source code in
-- return for reimbursement of the cost of distribution. This written offer
-- must permit verbatim duplication by anyone, or (C) it is distributed by
-- someone who received only the executable form, and is accompanied by a
-- copy of the written offer of source code.

-- 6. r-VEX was developed by Stephan Wong, Thijs van As, Fakhar Anjam,
-- Roel Seedorf, Anthony Brandon, Jeroen van Straten. r-VEX is currently
-- maintained by TU Delft (J.S.S.M.Wong@tudelft.nl).

-- 7. The MMU was developed by Jens Johansen.

-- Copyright (C) 2008-2016 by TU Delft.

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;


entity mmu_oh2bin is
  generic(
    WIDTH_LOG2                  : integer
  );
  port(
    oh_in                       : in  std_logic_vector(2**WIDTH_LOG2-1 downto 0);
    bin_out                     : out integer range 0 to 2**WIDTH_LOG2-1;
    hit                         : out std_logic
  );
end entity;

architecture log of mmu_oh2bin is 
  type t_valid_tree    is array (0 to WIDTH_LOG2-1)        of std_logic_vector(2**(WIDTH_LOG2 - 1) - 1 downto 0);
  type t_encode_vector is array (0 to 2**(WIDTH_LOG2-1)-1) of std_logic_vector(WIDTH_LOG2-1 downto 0);
  type t_encode_tree   is array (0 to WIDTH_LOG2-1)        of t_encode_vector;

  signal valid_tree  : t_valid_tree;
  signal encode_tree : t_encode_tree;

begin

  decoder_tree: process(oh_in, valid_tree, encode_tree) 
  begin 

    for lvl in 0 to WIDTH_LOG2-1 loop
      for i in 0 to 2**(WIDTH_LOG2-1-lvl) - 1 loop

        if lvl = 0 then
          valid_tree(0)(i)  <= oh_in(2 * i) or oh_in(2 * i + 1);
          encode_tree(0)(i)(0) <= oh_in(2 * i + 1);
        end if;

        if lvl > 0 then
          valid_tree(lvl)(i)  <= valid_tree(lvl - 1)(2 * i) or valid_tree(lvl - 1)(2 * i + 1);
        
          encode_tree(lvl)(i)(lvl) <= valid_tree(lvl - 1)(2 * i + 1);

          if valid_tree(lvl - 1)(2 * i + 1) = '1' then
            encode_tree(lvl)(i)(lvl-1 downto 0) <= encode_tree(lvl-1)(2 * i + 1)(lvl-1 downto 0);
          else
            encode_tree(lvl)(i)(lvl-1 downto 0) <= encode_tree(lvl-1)(2 * i)(lvl-1 downto 0);
          end if;
        end if;

      end loop;
    end loop;

  end process;

  hit   <= valid_tree(WIDTH_LOG2-1)(0);
  bin_out <= to_integer(unsigned(encode_tree(WIDTH_LOG2-1)(0)));

end architecture;