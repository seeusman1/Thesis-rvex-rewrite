-- Insert license here

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library work;
use work.rvex_pkg.all;
use work.rvex_intIface_pkg.all;

--=============================================================================
-- Testbench for the configuration control unit. It will attempt
-- reconfiguration to every runtime configuration which should be possible,
-- given a constant design time configuration. Conformance must be determined
-- manually from the simulation result for all design-time configurations.
-------------------------------------------------------------------------------
entity rvex_cfgCtrl_tb is
end rvex_cfgCtrl_tb;
--=============================================================================

--=============================================================================
architecture Behavioral of rvex_cfgCtrl_tb is
--=============================================================================
  
  -- rvex generic configuration.
  constant CFG                  : rvex_generic_config_type := (
    numLanesLog2                => 3,
    numLaneGroupsLog2           => 2,
    numContextsLog2             => 2,
    genBundleSizeLog2           => 3,
    multiplierLanes             => 2#11111111#,
    memLaneRevIndex             => 1,
    branchLaneRevIndex          => 0,
    numBreakpoints              => 4,
    forwarding                  => true,
    limmhFromNeighbor           => true,
    limmhFromPreviousPair       => true,
    reg63isLink                 => false,
    cregStartAddress            => X"FFFFFF80",
    resetVectors                => (others => (others => '0'))
  );
  
  -- Signals from and to the configuration controller.
  signal reset                       : std_logic;
  signal clk                         : std_logic;
  signal clkEn                       : std_logic;
  signal cxreg2cfg_requestData_r     : rvex_data_array(2**CFG.numContextsLog2-1 downto 0);
  signal cxreg2cfg_requestEnable     : std_logic_vector(2**CFG.numContextsLog2-1 downto 0);
  signal gbreg2cfg_requestData_r     : rvex_data_type;
  signal gbreg2cfg_requestEnable     : std_logic;
  signal cfg2gbreg_currentCfg        : rvex_data_type;
  signal cfg2gbreg_busy              : std_logic;
  signal cfg2gbreg_error             : std_logic;
  signal cfg2gbreg_requesterID       : std_logic_vector(3 downto 0);
  signal cfg2cxplif_run              : std_logic_vector(2**CFG.numContextsLog2-1 downto 0);
  signal cxplif2cfg_blockReconfig    : std_logic_vector(2**CFG.numContextsLog2-1 downto 0);
  signal mem2cfg_blockReconfig       : std_logic_vector(2**CFG.numLaneGroupsLog2-1 downto 0);
  signal cfg2any_coupled             : std_logic_vector(4**CFG.numLaneGroupsLog2-1 downto 0);
  signal cfg2any_decouple            : std_logic_vector(2**CFG.numLaneGroupsLog2-1 downto 0);
  signal cfg2any_numGroupsLog2       : rvex_2bit_array(2**CFG.numLaneGroupsLog2-1 downto 0);
  signal cfg2any_context             : rvex_3bit_array(2**CFG.numLaneGroupsLog2-1 downto 0);
  signal cfg2any_lastGroupForCtxt    : rvex_3bit_array(2**CFG.numContextsLog2-1 downto 0);
    
  -- Synchronization signal. This has a rising edge at every 10ns mark. It is
  -- used to align things to make them look nice in simulation.
  signal sync                        : std_logic := '0';
  
  -- Counts the number of valid configurations.
  signal validConfigs                : unsigned(31 downto 0);
  
--=============================================================================
begin
--=============================================================================
  
  -- Instantiate the configuration controller.
  uut: entity work.rvex_cfgCtrl
    generic map (
      CFG => CFG
    )
    port map (
      reset                       => reset,
      clk                         => clk,
      clkEn                       => clkEn,
      cxreg2cfg_requestData_r     => cxreg2cfg_requestData_r,
      cxreg2cfg_requestEnable     => cxreg2cfg_requestEnable,
      gbreg2cfg_requestData_r     => gbreg2cfg_requestData_r,
      gbreg2cfg_requestEnable     => gbreg2cfg_requestEnable,
      cfg2gbreg_currentCfg        => cfg2gbreg_currentCfg,
      cfg2gbreg_busy              => cfg2gbreg_busy,
      cfg2gbreg_error             => cfg2gbreg_error,
      cfg2gbreg_requesterID       => cfg2gbreg_requesterID,
      cfg2cxplif_run              => cfg2cxplif_run,
      cxplif2cfg_blockReconfig    => cxplif2cfg_blockReconfig,
      mem2cfg_blockReconfig       => mem2cfg_blockReconfig,
      cfg2any_coupled             => cfg2any_coupled,
      cfg2any_decouple            => cfg2any_decouple,
      cfg2any_numGroupsLog2       => cfg2any_numGroupsLog2,
      cfg2any_context             => cfg2any_context,
      cfg2any_lastGroupForCtxt    => cfg2any_lastGroupForCtxt
    );
  
  -- Drive the configuration block signals low, so reconfiguration is instant.
  cxplif2cfg_blockReconfig <= (others => '0');
  mem2cfg_blockReconfig <= (others => '0');
  
  -- Load default values into the requests from the contexts, we're not using
  -- them in this testbench.
  cxreg2cfg_requestData_r <= (others => (others => '0'));
  cxreg2cfg_requestEnable <= (others => '0');
  
  -- Generate sync signal.
  process is
  begin
    wait for 1 ps;
    sync <= '0';
    wait for 99999 ps;
    sync <= '1';
  end process;
  
  -- Generate other stimuli.
  process is
    type natural_array is array (natural range <>) of natural;
    variable contexts: natural_array(2**CFG.numLaneGroupsLog2-1 downto 0);
    variable carry: boolean;
    variable word: rvex_data_type;
  begin
    
    -- Reset everything.
    validConfigs <= (others => '0');
    gbreg2cfg_requestData_r <= (others => '0');
    gbreg2cfg_requestEnable <= '0';
    reset <= '1';
    clkEn <= '1';
    clk <= '1';
    wait for 1 ps;
    clk <= '0';
    wait for 1 ps;
    clk <= '1';
    wait for 1 ps;
    clk <= '0';
    wait for 1 ps;
    reset <= '0';
    
    -- Start out with everything connected to context 0.
    contexts := (others => 0);
    
    -- Loop over all configurations possible for 4-way reconfiguration, barring
    -- reserved bits.
    loop
      
      -- Encode the configuration word.
      word := (others => '0');
      for i in 0 to 2**CFG.numLaneGroupsLog2-1 loop
        if contexts(i) = 2**CFG.numContextsLog2 then
          
          -- Disable lane group.
          word(i*4+3) := '1';
          
        else
          
          -- Connect lane group to given context.
          word(i*4+CFG.numContextsLog2-1 downto i*4) :=
            std_logic_vector(to_unsigned(contexts(i), CFG.numContextsLog2));
          
        end if;
      end loop;
      
      -- Clock in the request.
      gbreg2cfg_requestEnable <= '1';
      wait for 1 ps;
      clk <= '1';
      wait for 1 ps;
      clk <= '0';
      gbreg2cfg_requestEnable <= '0';
      gbreg2cfg_requestData_r <= word;
      
      -- Send 10 clock pulses, after which reconfiguration should be complete.
      for i in 1 to 10 loop
        wait for 1 ps;
        clk <= '1';
        wait for 1 ps;
        clk <= '0';
      end loop;
      
      -- If the error bit is not set, this was considered to be a valid
      -- configuration. In that case, synchronize with the sync signal so the
      -- valid configuration words and their output can be easily seen.
      if cfg2gbreg_error = '0' then
        validConfigs <= validConfigs + 1;
        wait until rising_edge(sync);
      end if;
      
      -- Determine the next configuration to try.
      carry := true;
      for i in 0 to 2**CFG.numLaneGroupsLog2-1 loop
        contexts(i) := contexts(i) + 1;
        if contexts(i) = 2**CFG.numContextsLog2+1 then
          contexts(i) := 0;
        else
          carry := false;
          exit;
        end if;
      end loop;
      exit when carry;
      
    end loop;
    
    -- Stop simulation.
    report "Done!" severity failure;
    wait;
    
  end process;
  
end Behavioral;

