../../lib/rvex/core/core_opcode_pkg.template.vhd