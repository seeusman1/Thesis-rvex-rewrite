../../platform/core-tests/share/core_tb.template.vhd