../../lib/rvex/core/core_contextRegLogic.template.vhd