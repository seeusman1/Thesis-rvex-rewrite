-- r-VEX processor
-- Copyright (C) 2008-2016 by TU Delft.
-- All Rights Reserved.

-- THIS IS A LEGAL DOCUMENT, BY USING r-VEX,
-- YOU ARE AGREEING TO THESE TERMS AND CONDITIONS.

-- No portion of this work may be used by any commercial entity, or for any
-- commercial purpose, without the prior, written permission of TU Delft.
-- Nonprofit and noncommercial use is permitted as described below.

-- 1. r-VEX is provided AS IS, with no warranty of any kind, express
-- or implied. The user of the code accepts full responsibility for the
-- application of the code and the use of any results.

-- 2. Nonprofit and noncommercial use is encouraged. r-VEX may be
-- downloaded, compiled, synthesized, copied, and modified solely for nonprofit,
-- educational, noncommercial research, and noncommercial scholarship
-- purposes provided that this notice in its entirety accompanies all copies.
-- Copies of the modified software can be delivered to persons who use it
-- solely for nonprofit, educational, noncommercial research, and
-- noncommercial scholarship purposes provided that this notice in its
-- entirety accompanies all copies.

-- 3. ALL COMMERCIAL USE, AND ALL USE BY FOR PROFIT ENTITIES, IS EXPRESSLY
-- PROHIBITED WITHOUT A LICENSE FROM TU Delft (J.S.S.M.Wong@tudelft.nl).

-- 4. No nonprofit user may place any restrictions on the use of this software,
-- including as modified by the user, by any other authorized user.

-- 5. Noncommercial and nonprofit users may distribute copies of r-VEX
-- in compiled or binary form as set forth in Section 2, provided that
-- either: (A) it is accompanied by the corresponding machine-readable source
-- code, or (B) it is accompanied by a written offer, with no time limit, to
-- give anyone a machine-readable copy of the corresponding source code in
-- return for reimbursement of the cost of distribution. This written offer
-- must permit verbatim duplication by anyone, or (C) it is distributed by
-- someone who received only the executable form, and is accompanied by a
-- copy of the written offer of source code.

-- 6. r-VEX was developed by Stephan Wong, Thijs van As, Fakhar Anjam,
-- Roel Seedorf, Anthony Brandon, Jeroen van Straten. r-VEX is currently
-- maintained by TU Delft (J.S.S.M.Wong@tudelft.nl).

-- Copyright (C) 2008-2016 by TU Delft.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library rvex;
use rvex.common_pkg.all;
use rvex.utils_pkg.all;
use rvex.cache_pkg.all;

entity cache_tlb_cams_tb is
end cache_tlb_cams_tb;

architecture testbench of cache_tlb_cams_tb is
  
  -- UUT generics.
  constant CCFG : cache_generic_config_type := cache_cfg(
    camStyle => CRS_BRAM36
  );
  
  -- UUT signals.
  signal reset                  : std_logic;
  signal resetting              : std_logic;
  signal clk                    : std_logic;
  signal vAddr                  : rvex_address_type;
  signal asid                   : rvex_data_type;
  signal entry_valid            : std_logic;
  signal entry_index            : std_logic_vector(CCFG.tlbDepthLog2-1 downto 0);
  signal entry_global           : std_logic;
  signal entry_large            : std_logic;
  signal update_op              : std_logic_vector(1 downto 0);
  signal update_index           : std_logic_vector(CCFG.tlbDepthLog2-1 downto 0);
  signal update_global          : std_logic;
  signal update_large           : std_logic;
  
begin
  
  -- Instantiate UUT.
  uut: entity work.cache_tlb_cams
    generic map (
      CCFG          => CCFG
    )
    port map (
      
      -- System control.
      reset         => reset,
      resetting     => resetting,
      clk           => clk,
      
      -- CAM read port.
      vAddr         => vAddr,
      asid          => asid,
      entry_valid   => entry_valid,
      entry_index   => entry_index,
      entry_global  => entry_global,
      entry_large   => entry_large,
      
      -- CAM write port.
      update_op     => update_op,
      update_index  => update_index,
      update_global => update_global,
      update_large  => update_large
      
    );
  
  -- Generate clock.
  clk_proc: process is
  begin
    clk <= '1';
    wait for 5 ns;
    clk <= '0';
    wait for 5 ns;
  end process;
  
  -- Generate stimuli.
  stim_proc: process is
  begin
    
    -- Assign undefined to all inputs except for the command input, which we
    -- assign to no-operation.
    vAddr         <= (others => 'U');
    asid          <= (others => 'U');
    update_op     <= "00";
    update_index  <= (others => 'U');
    update_global <= 'U';
    update_large  <= 'U';
    
    -- Assert reset for two cycles.
    reset <= '1';
    wait until rising_edge(clk);
    wait until rising_edge(clk);
    reset <= '0';
    
    -- Wait until the CAM finishes resetting.
    wait until rising_edge(clk) and resetting = '0';
    
    wait;
  end process;
  
end testbench;

