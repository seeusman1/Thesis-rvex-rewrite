-- r-VEX processor
-- Copyright (C) 2008-2014 by TU Delft.
-- All Rights Reserved.

-- THIS IS A LEGAL DOCUMENT, BY USING r-VEX,
-- YOU ARE AGREEING TO THESE TERMS AND CONDITIONS.

-- No portion of this work may be used by any commercial entity, or for any
-- commercial purpose, without the prior, written permission of TU Delft.
-- Nonprofit and noncommercial use is permitted as described below.

-- 1. r-VEX is provided AS IS, with no warranty of any kind, express
-- or implied. The user of the code accepts full responsibility for the
-- application of the code and the use of any results.

-- 2. Nonprofit and noncommercial use is encouraged. r-VEX may be
-- downloaded, compiled, synthesized, copied, and modified solely for nonprofit,
-- educational, noncommercial research, and noncommercial scholarship
-- purposes provided that this notice in its entirety accompanies all copies.
-- Copies of the modified software can be delivered to persons who use it
-- solely for nonprofit, educational, noncommercial research, and
-- noncommercial scholarship purposes provided that this notice in its
-- entirety accompanies all copies.

-- 3. ALL COMMERCIAL USE, AND ALL USE BY FOR PROFIT ENTITIES, IS EXPRESSLY
-- PROHIBITED WITHOUT A LICENSE FROM TU Delft (J.S.S.M.Wong@tudelft.nl).

-- 4. No nonprofit user may place any restrictions on the use of this software,
-- including as modified by the user, by any other authorized user.

-- 5. Noncommercial and nonprofit users may distribute copies of r-VEX
-- in compiled or binary form as set forth in Section 2, provided that
-- either: (A) it is accompanied by the corresponding machine-readable source
-- code, or (B) it is accompanied by a written offer, with no time limit, to
-- give anyone a machine-readable copy of the corresponding source code in
-- return for reimbursement of the cost of distribution. This written offer
-- must permit verbatim duplication by anyone, or (C) it is distributed by
-- someone who received only the executable form, and is accompanied by a
-- copy of the written offer of source code.

-- 6. r-VEX was developed by Stephan Wong, Thijs van As, Fakhar Anjam,
-- Roel Seedorf, Anthony Brandon, Jeroen van Straten. r-VEX is currently
-- maintained by TU Delft (J.S.S.M.Wong@tudelft.nl).

-- Copyright (C) 2008-2014 by TU Delft.

-- Refer to reconfCache_pkg.vhd for configuration constants and most
-- documentation.

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library rvex;
use rvex.cache_pkg.all;

entity cache_tb_mockMemBus is
  port (
    
    -- Clock input.
    clk                       : in  std_logic;
    
    -- Active high reset input.
    reset                     : in  std_logic;
    
    -- Active high clock enable input.
    clkEn                     : in  std_logic;
    
    -- Bus masters.
    arbToCache                : out reconfCache_memIn_array;
    cacheToArb                : in  reconfCache_memOut_array;
    
    -- Arbitrated bus output.
    memToArb                  : in  reconfCache_memIn;
    arbToMem                  : out reconfCache_memOut
    
  );
end cache_tb_mockMemBus;

architecture Behavioral of cache_tb_mockMemBus is
  
  -- State machine state/mux selection signals.
  signal selectCache_next     : natural;
  signal selectCache          : natural;
  
begin
  
  --===========================================================================
  -- Generate mux/demux logic
  --===========================================================================
  to_masters_gen: for i in 0 to RC_NUM_ATOMS-1 generate
    arbToCache(i).ready <= memToArb.ready when selectCache = i else '0';
    arbToCache(i).data  <= memToArb.data;
  end generate;
  
  arbToMem.addr         <= cacheToArb(selectCache_next).addr;
  arbToMem.readEnable   <= cacheToArb(selectCache_next).readEnable;
  arbToMem.writeData    <= cacheToArb(selectCache_next).writeData;
  arbToMem.writeMask    <= cacheToArb(selectCache_next).writeMask;
  arbToMem.writeEnable  <= cacheToArb(selectCache_next).writeEnable;
  arbToMem.burstEnable  <= cacheToArb(selectCache_next).burstEnable;
  
  --===========================================================================
  -- Generate the selection state machine
  --===========================================================================
  select_comb: process (memToArb.ready, selectCache, cacheToArb) is
  begin
    if memToArb.ready = '1' then
      
      -- If the currently selected master is not accessing the bus, move to the
      -- next.
      if cacheToArb(selectCache).readEnable = '0' and cacheToArb(selectCache).writeEnable = '0' then
        if selectCache >= RC_NUM_ATOMS-1 then
          selectCache_next <= 0;
        else
          selectCache_next <= selectCache + 1;
        end if;
      end if;
      
    else
      
      -- Switching is not allowed in the middle of a transaction.
      selectCache_next <= selectCache;
      
    end if;
  end process;
  
  select_seq: process (clk) is
  begin
    if rising_edge(clk) then
      if reset = '1' then
        selectCache <= 0;
      elsif clkEn = '1' then
        selectCache <= selectCache_next;
      end if;
    end if;
  end process;
  
end Behavioral;

